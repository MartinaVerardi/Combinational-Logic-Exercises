/*

A) Write a systemVerilog module that calculates the day of the year, e.g., 
February 1 would be the day 32nd day of the year. Ignore leap years for now. 
The header for the module is:

module dayIfYrCalc
    (
    input logic [5:0] dayOfMonth,
    input logic [3:0] month,
    output logic [8:0] dayOfYear;
    );

*/